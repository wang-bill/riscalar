fjkdsa
