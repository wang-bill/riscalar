`timescale 1ns / 1ps
`default_nettype none

module register_file
  (
    input wire [4:0] rs1_in,
    input wire [4:0] rs2_in,
    
  )

endmodule

`default_nettype wire